* T29U SPICE BSIM3 VERSION 3.1 PARAMETERS

*SPICE 3f5 Level 8, Star-HSPICE Level 49, UTMOST Level 8

* DATE: Nov  6/02
* LOT: T29U                  WAF: 8001
* Temperature_parameters=Default
.MODEL NMOS NMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 5.7E-9
+XJ      = 1E-7           NCH     = 2.3549E17      VTH0    = 0.388582
+K1      = 0.4545906      K2      = 4.630687E-3    K3      = 1E-3
+K3B     = 2.7003371      W0      = 1E-7           NLX     = 2.469653E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 0.360271       DVT1    = 0.3829891      DVT2    = -0.5
+U0      = 304.6846051    UA      = -1.174063E-9   UB      = 2.397658E-18
+UC      = 3.541076E-11   VSAT    = 1.539191E5     A0      = 1.6070193
+AGS     = 0.2905776      B0      = -1.854529E-7   B1      = 8.598488E-7
+KETA    = -1.783772E-3   A1      = 1.916643E-4    A2      = 0.4162048
+RDSW    = 133.8002918    PRWG    = 0.5            PRWB    = -0.2
+WR      = 1              WINT    = 0              LINT    = 8.641225E-9
+XL      = 3E-8           XW      = -4E-8          DWG     = -1.189337E-8
+DWB     = 4.492511E-9    VOFF    = -0.0984831     NFACTOR = 1.8462358
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 5.063972E-3    ETAB    = 5.522478E-4
+DSUB    = 0.0306469      PCLM    = 1.801348       PDIBLC1 = 1
+PDIBLC2 = 2.698952E-3    PDIBLCB = -0.0911843     DROUT   = 0.9029812
+PSCBE1  = 7.995457E10    PSCBE2  = 5.012176E-10   PVAG    = 0
+DELTA   = 0.01           RSH     = 4.7            MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 5.7E-10        CGSO    = 5.7E-10        CGBO    = 1E-12
+CJ      = 1.692268E-3    PB      = 0.99           MJ      = 0.4461196
+CJSW    = 3.80197E-10    PBSW    = 0.860409       MJSW    = 0.3703426
+CJSWG   = 3.29E-10       PBSWG   = 0.860409       MJSWG   = 0.3703426
+CF      = 0              PVTH0   = -8.610903E-3   PRDSW   = -10
+PK2     = 3.16474E-3     WKETA   = 3.726252E-3    LKETA   = -8.399886E-3    )
*
.MODEL PMOS PMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 5.7E-9
+XJ      = 1E-7           NCH     = 4.1589E17      VTH0    = -0.5538459
+K1      = 0.6241479      K2      = 1.799564E-3    K3      = 0
+K3B     = 12.9869461     W0      = 1E-6           NLX     = 1E-9
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 3.4046733      DVT1    = 0.8388132      DVT2    = -0.1233861
+U0      = 108.1056054    UA      = 1.268292E-9    UB      = 1.168491E-21
+UC      = -1E-10         VSAT    = 2E5            A0      = 0.9429827
+AGS     = 0.1779362      B0      = 1.186871E-6    B1      = 5E-6
+KETA    = 0.0181651      A1      = 6.003832E-3    A2      = 0.3
+RDSW    = 769.9250696    PRWG    = 0.3542925      PRWB    = -0.3256606
+WR      = 1              WINT    = 0              LINT    = 4.151327E-8
+XL      = 3E-8           XW      = -4E-8          DWG     = -3.684793E-8
+DWB     = 6.196368E-9    VOFF    = -0.1316705     NFACTOR = 1.045776
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 0.5610656      ETAB    = -0.0743897
+DSUB    = 1.1987358      PCLM    = 1.254027       PDIBLC1 = 5.616609E-3
+PDIBLC2 = 9.953866E-9    PDIBLCB = -6.082702E-4   DROUT   = 0.0786297
+PSCBE1  = 3.266969E9     PSCBE2  = 6.01449E-10    PVAG    = 8.90109E-3
+DELTA   = 0.01           RSH     = 3.5            MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 6.6E-10        CGSO    = 6.6E-10        CGBO    = 1E-12
+CJ      = 1.896791E-3    PB      = 0.99           MJ      = 0.4683049
+CJSW    = 3.502714E-10   PBSW    = 0.6971859      MJSW    = 0.2558685
+CJSWG   = 2.5E-10        PBSWG   = 0.6971859      MJSWG   = 0.2558685
+CF      = 0              PVTH0   = 4.759823E-3    PRDSW   = 10.0559187
+PK2     = 2.906223E-3    WKETA   = 0.0252043      LKETA   = -0.010831       )
*